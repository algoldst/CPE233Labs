`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly
// Engineer: Paul Hummel
//
// Create Date: 06/28/2018 05:21:01 AM
// Module Name: RAT_WRAPPER
// Target Devices: RAT MCU on Basys3
// Description: Basic RAT_WRAPPER
//
// Revision:
// Revision 0.01 - File Created
//////////////////////////////////////////////////////////////////////////////

module Rat_Wrapper(
    input CLK,
    input BTNC,
    input BTNL,
    input [7:0] SWITCHES,
    output [7:0] LEDS,
    output [7:0] SSEG, // SSEG segments
    output [3:0] DISP_EN // SSEG on/off
    );
    
    // INPUT PORT IDS ////////////////////////////////////////////////////////
    // Right now, the only possible inputs are the switches
    // In future labs you can add more port IDs, and you'll have
    // to add constants here for the mux below
    localparam SWITCHES_ID = 8'h20;
       
    // OUTPUT PORT IDS ///////////////////////////////////////////////////////
    // In future labs you can add more port IDs
    localparam LEDS_ID      = 8'h40;
    localparam SSEG_ID      = 8'h81;
       
    // Signals for connecting RAT_MCU to RAT_wrapper /////////////////////////
    logic [7:0] s_output_port;
    logic [7:0] s_port_id;
    logic s_load;
    logic s_interrupt;
    logic s_reset;
    logic s_clk_50 = 1'b0;     // 50 MHz clock
    logic btn_debounce;
    
    // Register definitions for output devices ///////////////////////////////
    logic [7:0]   s_input_port;
    logic [7:0]   r_leds = 8'h00;
    logic [15:0]   r_sseg = 8'h00;

    // Declare RAT_CPU ///////////////////////////////////////////////////////
    MCU MCU(.in_port(s_input_port), .out_port(s_output_port),
                .port_id(s_port_id), .io_strb(s_load), .reset(s_reset),
                .interrupt(s_interrupt /*BTNL*/), .clk(s_clk_50)); //BTNL for bypassing Debounce (do this in Sim!)
    
    // Clock Divider to create 50 MHz Clock //////////////////////////////////
    always_ff @(posedge CLK) begin
        s_clk_50 <= ~s_clk_50;
    end
    
     
    // MUX for selecting what input to read //////////////////////////////////
    always_comb begin
        if (s_port_id == SWITCHES_ID)
            s_input_port = SWITCHES;
        else
            s_input_port = 8'h00;
    end
   
    // MUX for updating output registers /////////////////////////////////////
    // Register updates depend on rising clock edge and asserted load signal
    always_ff @ (posedge CLK) begin
        if (s_load == 1'b1) begin
            if (s_port_id == LEDS_ID)
                r_leds <= s_output_port;
            else if (s_port_id == SSEG_ID)
                r_sseg <= s_output_port;
        end
    end
     
    // Connect Signals ///////////////////////////////////////////////////////
    assign s_reset = BTNC;
    //assign s_interrupt = 1'b0;  // no interrupt used yet
     
    // Output Assignments ////////////////////////////////////////////////////
    assign LEDS = r_leds;
   
    // SSEG Display    ////////////////////////////////////////////////////
    SevSegDisp sseg(.CLK(CLK), .MODE(0), .DATA_IN(r_sseg), .CATHODES(SSEG), 
                    .ANODES(DISP_EN) );  
   // Debounce Circuit
    Debounce debounce(.CLK(CLK), .BTN(BTNL), .DB_BTN(s_interrupt));
    endmodule
